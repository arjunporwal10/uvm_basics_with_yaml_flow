`ifndef EXAMPLE_BUS_SEQ_LIST__SV
`define EXAMPLE_BUS_SEQ_LIST__SV

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "example_bus_write_seq.sv"
`include "example_bus_read_seq.sv"

`endif
